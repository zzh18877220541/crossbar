module crossbar64x64 #(
    parameter width = 320,
    parameter depth1 = 64,
    parameter depth2 = 128,
)(
    input wire [5:0] sel_in0,
    input wire [width - 1:0] in0,
    input wire [5:0] sel_in1,
    input wire [width - 1:0] in1,
    input wire [5:0] sel_in2,
    input wire [width - 1:0] in2,
    input wire [5:0] sel_in3,
    input wire [width - 1:0] in3,
    input wire [5:0] sel_in4,
    input wire [width - 1:0] in4,
    input wire [5:0] sel_in5,
    input wire [width - 1:0] in5,
    input wire [5:0] sel_in6,
    input wire [width - 1:0] in6,
    input wire [5:0] sel_in7,
    input wire [width - 1:0] in7,
    input wire [5:0] sel_in8,
    input wire [width - 1:0] in8,
    input wire [5:0] sel_in9,
    input wire [width - 1:0] in9,
    input wire [5:0] sel_in10,
    input wire [width - 1:0] in10,
    input wire [5:0] sel_in11,
    input wire [width - 1:0] in11,
    input wire [5:0] sel_in12,
    input wire [width - 1:0] in12,
    input wire [5:0] sel_in13,
    input wire [width - 1:0] in13,
    input wire [5:0] sel_in14,
    input wire [width - 1:0] in14,
    input wire [5:0] sel_in15,
    input wire [width - 1:0] in15,
    input wire [5:0] sel_in16,
    input wire [width - 1:0] in16,
    input wire [5:0] sel_in17,
    input wire [width - 1:0] in17,
    input wire [5:0] sel_in18,
    input wire [width - 1:0] in18,
    input wire [5:0] sel_in19,
    input wire [width - 1:0] in19,
    input wire [5:0] sel_in20,
    input wire [width - 1:0] in20,
    input wire [5:0] sel_in21,
    input wire [width - 1:0] in21,
    input wire [5:0] sel_in22,
    input wire [width - 1:0] in22,
    input wire [5:0] sel_in23,
    input wire [width - 1:0] in23,
    input wire [5:0] sel_in24,
    input wire [width - 1:0] in24,
    input wire [5:0] sel_in25,
    input wire [width - 1:0] in25,
    input wire [5:0] sel_in26,
    input wire [width - 1:0] in26,
    input wire [5:0] sel_in27,
    input wire [width - 1:0] in27,
    input wire [5:0] sel_in28,
    input wire [width - 1:0] in28,
    input wire [5:0] sel_in29,
    input wire [width - 1:0] in29,
    input wire [5:0] sel_in30,
    input wire [width - 1:0] in30,
    input wire [5:0] sel_in31,
    input wire [width - 1:0] in31,
    input wire [5:0] sel_in32,
    input wire [width - 1:0] in32,
    input wire [5:0] sel_in33,
    input wire [width - 1:0] in33,
    input wire [5:0] sel_in34,
    input wire [width - 1:0] in34,
    input wire [5:0] sel_in35,
    input wire [width - 1:0] in35,
    input wire [5:0] sel_in36,
    input wire [width - 1:0] in36,
    input wire [5:0] sel_in37,
    input wire [width - 1:0] in37,
    input wire [5:0] sel_in38,
    input wire [width - 1:0] in38,
    input wire [5:0] sel_in39,
    input wire [width - 1:0] in39,
    input wire [5:0] sel_in40,
    input wire [width - 1:0] in40,
    input wire [5:0] sel_in41,
    input wire [width - 1:0] in41,
    input wire [5:0] sel_in42,
    input wire [width - 1:0] in42,
    input wire [5:0] sel_in43,
    input wire [width - 1:0] in43,
    input wire [5:0] sel_in44,
    input wire [width - 1:0] in44,
    input wire [5:0] sel_in45,
    input wire [width - 1:0] in45,
    input wire [5:0] sel_in46,
    input wire [width - 1:0] in46,
    input wire [5:0] sel_in47,
    input wire [width - 1:0] in47,
    input wire [5:0] sel_in48,
    input wire [width - 1:0] in48,
    input wire [5:0] sel_in49,
    input wire [width - 1:0] in49,
    input wire [5:0] sel_in50,
    input wire [width - 1:0] in50,
    input wire [5:0] sel_in51,
    input wire [width - 1:0] in51,
    input wire [5:0] sel_in52,
    input wire [width - 1:0] in52,
    input wire [5:0] sel_in53,
    input wire [width - 1:0] in53,
    input wire [5:0] sel_in54,
    input wire [width - 1:0] in54,
    input wire [5:0] sel_in55,
    input wire [width - 1:0] in55,
    input wire [5:0] sel_in56,
    input wire [width - 1:0] in56,
    input wire [5:0] sel_in57,
    input wire [width - 1:0] in57,
    input wire [5:0] sel_in58,
    input wire [width - 1:0] in58,
    input wire [5:0] sel_in59,
    input wire [width - 1:0] in59,
    input wire [5:0] sel_in60,
    input wire [width - 1:0] in60,
    input wire [5:0] sel_in61,
    input wire [width - 1:0] in61,
    input wire [5:0] sel_in62,
    input wire [width - 1:0] in62,
    input wire [5:0] sel_in63,
    input wire [width - 1:0] in63,
    input wire clk,
    input wire rst,
    output reg [width - 1:0] out0,
    output reg [width - 1:0] out1,
    output reg [width - 1:0] out2,
    output reg [width - 1:0] out3,
    output reg [width - 1:0] out4,
    output reg [width - 1:0] out5,
    output reg [width - 1:0] out6,
    output reg [width - 1:0] out7,
    output reg [width - 1:0] out8,
    output reg [width - 1:0] out9,
    output reg [width - 1:0] out10,
    output reg [width - 1:0] out11,
    output reg [width - 1:0] out12,
    output reg [width - 1:0] out13,
    output reg [width - 1:0] out14,
    output reg [width - 1:0] out15,
    output reg [width - 1:0] out16,
    output reg [width - 1:0] out17,
    output reg [width - 1:0] out18,
    output reg [width - 1:0] out19,
    output reg [width - 1:0] out20,
    output reg [width - 1:0] out21,
    output reg [width - 1:0] out22,
    output reg [width - 1:0] out23,
    output reg [width - 1:0] out24,
    output reg [width - 1:0] out25,
    output reg [width - 1:0] out26,
    output reg [width - 1:0] out27,
    output reg [width - 1:0] out28,
    output reg [width - 1:0] out29,
    output reg [width - 1:0] out30,
    output reg [width - 1:0] out31,
    output reg [width - 1:0] out32,
    output reg [width - 1:0] out33,
    output reg [width - 1:0] out34,
    output reg [width - 1:0] out35,
    output reg [width - 1:0] out36,
    output reg [width - 1:0] out37,
    output reg [width - 1:0] out38,
    output reg [width - 1:0] out39,
    output reg [width - 1:0] out40,
    output reg [width - 1:0] out41,
    output reg [width - 1:0] out42,
    output reg [width - 1:0] out43,
    output reg [width - 1:0] out44,
    output reg [width - 1:0] out45,
    output reg [width - 1:0] out46,
    output reg [width - 1:0] out47,
    output reg [width - 1:0] out48,
    output reg [width - 1:0] out49,
    output reg [width - 1:0] out50,
    output reg [width - 1:0] out51,
    output reg [width - 1:0] out52,
    output reg [width - 1:0] out53,
    output reg [width - 1:0] out54,
    output reg [width - 1:0] out55,
    output reg [width - 1:0] out56,
    output reg [width - 1:0] out57,
    output reg [width - 1:0] out58,
    output reg [width - 1:0] out59,
    output reg [width - 1:0] out60,
    output reg [width - 1:0] out61,
    output reg [width - 1:0] out62,
    output reg [width - 1:0] out63
);

reg [width - 1: 0] Group[3: 0][15: 0];

// Inputs
wire [width - 1: 0] in[63: 0]; // 16 input ports
wire [5: 0] sel_in[63: 0];    // 16 select signals

// Outputs
wire [width-1:0] out[63:0]; // 16 output ports

assign in[0] = in0, in[1] = in1, in[2] = in2, in[3] = in3, in[4] = in4, in[5] = in5, in[6] = in6, in[7] = in7, in[8] = in8, in[9] = in9, 
    in[10] = in10, in[11] = in11, in[12] = in12, in[13] = in13, in[14] = in14, in[15] = in15, in[16] = in16, in[17] = in17, 
    in[18] = in18, in[19] = in19, in[20] = in20, in[21] = in21, in[22] = in22, in[23] = in23, in[24] = in24, in[25] = in25, 
    in[26] = in26, in[27] = in27, in[28] = in28, in[29] = in29, in[30] = in30, in[31] = in31, in[32] = in32, in[33] = in33, 
    in[34] = in34, in[35] = in35, in[36] = in36, in[37] = in37, in[38] = in38, in[39] = in39, in[40] = in40, in[41] = in41, 
    in[42] = in42, in[43] = in43, in[44] = in44, in[45] = in45, in[46] = in46, in[47] = in47, in[48] = in48, in[49] = in49, 
    in[50] = in50, in[51] = in51, in[52] = in52, in[53] = in53, in[54] = in54, in[55] = in55, in[56] = in56, in[57] = in57, 
    in[58] = in58, in[59] = in59, in[60] = in60, in[61] = in61, in[62] = in62, in[63] = in63;

assign sel_in[0] = sel_in0, sel_in[1] = sel_in1, sel_in[2] = sel_in2, sel_in[3] = sel_in3, sel_in[4] = sel_in4, sel_in[5] = sel_in5, 
    sel_in[6] = sel_in6, sel_in[7] = sel_in7, sel_in[8] = sel_in8, sel_in[9] = sel_in9, sel_in[10] = sel_in10, sel_in[11] = sel_in11, 
    sel_in[12] = sel_in12, sel_in[13] = sel_in13, sel_in[14] = sel_in14, sel_in[15] = sel_in15, sel_in[16] = sel_in16, sel_in[17] = sel_in17, 
    sel_in[18] = sel_in18, sel_in[19] = sel_in19, sel_in[20] = sel_in20, sel_in[21] = sel_in21, sel_in[22] = sel_in22, sel_in[23] = sel_in23, 
    sel_in[24] = sel_in24, sel_in[25] = sel_in25, sel_in[26] = sel_in26, sel_in[27] = sel_in27, sel_in[28] = sel_in28, sel_in[29] = sel_in29, 
    sel_in[30] = sel_in30, sel_in[31] = sel_in31, sel_in[32] = sel_in32, sel_in[33] = sel_in33, sel_in[34] = sel_in34, sel_in[35] = sel_in35, 
    sel_in[36] = sel_in36, sel_in[37] = sel_in37, sel_in[38] = sel_in38, sel_in[39] = sel_in39, sel_in[40] = sel_in40, sel_in[41] = sel_in41, 
    sel_in[42] = sel_in42, sel_in[43] = sel_in43, sel_in[44] = sel_in44, sel_in[45] = sel_in45, sel_in[46] = sel_in46, sel_in[47] = sel_in47, 
    sel_in[48] = sel_in48, sel_in[49] = sel_in49, sel_in[50] = sel_in50, sel_in[51] = sel_in51, sel_in[52] = sel_in52, sel_in[53] = sel_in53,
    sel_in[54] = sel_in54, sel_in[55] = sel_in55, sel_in[56] = sel_in56, sel_in[57] = sel_in57, sel_in[58] = sel_in58, sel_in[59] = sel_in59,
    sel_in[60] = sel_in60, sel_in[61] = sel_in61, sel_in[62] = sel_in62, sel_in[63] = sel_in63;

assign out0 = out[0], out1 = out[1], out2 = out[2], out3 = out[3], out4 = out[4], out5 = out[5], out6 = out[6], out7 = out[7], 
    out8 = out[8], out9 = out[9], out10 = out[10], out11 = out[11], out12 = out[12], out13 = out[13], out14 = out[14], out15 = out[15], 
    out16 = out[16], out17 = out[17], out18 = out[18], out19 = out[19], out20 = out[20], out21 = out[21], out22 = out[22], out23 = out[23], 
    out24 = out[24], out25 = out[25], out26 = out[26], out27 = out[27], out28 = out[28], out29 = out[29], out30 = out[30], out31 = out[31], 
    out32 = out[32], out33 = out[33], out34 = out[34], out35 = out[35], out36 = out[36], out37 = out[37], out38 = out[38], out39 = out[39], 
    out40 = out[40], out41 = out[41], out42 = out[42], out43 = out[43], out44 = out[44], out45 = out[45], out46 = out[46], out47 = out[47], 
    out48 = out[48], out49 = out[49], out50 = out[50], out51 = out[51], out52 = out[52], out53 = out[53], out54 = out[54], out55 = out[55], 
    out56 = out[56], out57 = out[57], out58 = out[58], out59 = out[59], out60 = out[60], out61 = out[61], out62 = out[62], out63 = out[63];

genvar i;

gennerate
    for (i = 0; i < 16; i = i + 1) begin: 4x4
        crossbar4x4 #(
            .width(width),
            .depth(depth1)
        ) crossbar4x4 (
            .sel_in0(sel_in[i * 4 + 0]),
            .in0(in[i * 4 + 0]),
            .sel_in1(sel_in[i * 4 + 1]),
            .in1(in[i * 4 + 1]),
            .sel_in2(sel_in[i * 4 + 2]),
            .in2(in[i * 4 + 2]),
            .sel_in3(sel_in[i * 4 + 3]),
            .in3(in[i * 4 + 3]),
            .out0(out[i * 4 + 0]),
            .out1(out[i * 4 + 1]),
            .out2(out[i * 4 + 2]),
            .out3(out[i * 4 + 3]),
            .clk(clk),
            .rst(rst)
        );
    end
endgennerate

gennerate
    for (i = 0; i < 4; i = i + 1) begin: 16x16
        crossbar16x16 #(
            .width(width),
            .depth(depth2)
        ) crossbar16x16 (
            in0(in[i * 16 + 0]),
            in1(in[i * 16 + 1]),
            in2(in[i * 16 + 2]),
            in3(in[i * 16 + 3]),
            in4(in[i * 16 + 4]),
            in5(in[i * 16 + 5]),
            in6(in[i * 16 + 6]),
            in7(in[i * 16 + 7]),
            in8(in[i * 16 + 8]),
            in9(in[i * 16 + 9]),
            in10(in[i * 16 + 10]),
            in11(in[i * 16 + 11]),
            in12(in[i * 16 + 12]),
            in13(in[i * 16 + 13]),
            in14(in[i * 16 + 14]),
            in15(in[i * 16 + 15]),
            out0(Group[i][0]),
            out1(Group[i][1]),
            out2(Group[i][2]),
            out3(Group[i][3]),
            out4(Group[i][4]),
            out5(Group[i][5]),
            out6(Group[i][6]),
            out7(Group[i][7]),
            out8(Group[i][8]),
            out9(Group[i][9]),
            out10(Group[i][10]),
            out11(Group[i][11]),
            out12(Group[i][12]),
            out13(Group[i][13]),
            out14(Group[i][14]),
            out15(Group[i][15]),
            sel_in0(sel_in[i * 16 + 0]),
            sel_in1(sel_in[i * 16 + 1]),
            sel_in2(sel_in[i * 16 + 2]),
            sel_in3(sel_in[i * 16 + 3]),
            sel_in4(sel_in[i * 16 + 4]),
            sel_in5(sel_in[i * 16 + 5]),
            sel_in6(sel_in[i * 16 + 6]),
            sel_in7(sel_in[i * 16 + 7]),
            sel_in8(sel_in[i * 16 + 8]),
            sel_in9(sel_in[i * 16 + 9]),
            sel_in10(sel_in[i * 16 + 10]),
            sel_in11(sel_in[i * 16 + 11]),
            sel_in12(sel_in[i * 16 + 12]),
            sel_in13(sel_in[i * 16 + 13]),
            sel_in14(sel_in[i * 16 + 14]),
            sel_in15(sel_in[i * 16 + 15]),
            clk(clk),
            rst(rst)
        );
    end
endgennerate

endmodule
